LIBRARY ieee ;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all;
package pacote is
	type char_array is array (39 downto 0) of std_logic_vector(1 downto 0);
end pacote;