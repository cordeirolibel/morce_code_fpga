LIBRARY ieee;
USE ieee.std_logic_1164.all;
	
package meupacote is
	type SSDARRAY is array (natural range <>) of STD_LOGIC_VECTOR (0 TO 6);
	
	CONSTANT num_0 : STD_LOGIC_VECTOR (0 TO 6) := "0000001";
	CONSTANT num_1 : STD_LOGIC_VECTOR (0 TO 6) := "1001111";
	CONSTANT num_2 : STD_LOGIC_VECTOR (0 TO 6) := "0010010";
	CONSTANT num_3 : STD_LOGIC_VECTOR (0 TO 6) := "0000110";
	CONSTANT num_4 : STD_LOGIC_VECTOR (0 TO 6) := "1001100";
	CONSTANT num_5 : STD_LOGIC_VECTOR (0 TO 6) := "0100100";
	CONSTANT num_6 : STD_LOGIC_VECTOR (0 TO 6) := "0100000";
	CONSTANT num_7 : STD_LOGIC_VECTOR (0 TO 6) := "0001111";
	CONSTANT num_8 : STD_LOGIC_VECTOR (0 TO 6) := "0000000";
	CONSTANT num_9 : STD_LOGIC_VECTOR (0 TO 6) := "0001100";
	CONSTANT num_a : STD_LOGIC_VECTOR (0 TO 6) := "0001000";
	CONSTANT num_b : STD_LOGIC_VECTOR (0 TO 6) := "1100000";
	CONSTANT num_c : STD_LOGIC_VECTOR (0 TO 6) := "0110001";
	CONSTANT num_d : STD_LOGIC_VECTOR (0 TO 6) := "1000010";
	CONSTANT num_e : STD_LOGIC_VECTOR (0 TO 6) := "0110000";
	CONSTANT num_f : STD_LOGIC_VECTOR (0 TO 6) := "0111000";
	CONSTANT negat : STD_LOGIC_VECTOR (0 TO 6) := "1111110";
	CONSTANT posit : STD_LOGIC_VECTOR (0 TO 6) := "1111111";
end package;