library ieee;

use ieee.std_logic_1164.all;

package mensagem is

--------------------------------------------------
TYPE char_array IS ARRAY (38 DOWNTO 0) OF std_logic_vector (1 DOWNTO 0); 
--------------------------------------------------


END mensagem;